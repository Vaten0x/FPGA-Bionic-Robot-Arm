module button_input(

);

endmodule;